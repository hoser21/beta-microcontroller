// ---------------------------------------------------------------------
//    Module:     32-bit CPU Data Path
//    Author:     Kevin Hoser and Alex Schendel
//    Contact:    hoser21@up.edu and schendel21@up.edu
//    Date:       5/11/2020
// ---------------------------------------------------------------------

`include "header.vh"

module CPUDataPath;